package spi_driver_pkg;

class spi_driver;



endclass

endpackage